`timescale 1ns / 1ps



module Extraction_Tb();

	reg [8:0]numberIn_tb;
	wire [6:0]whole;
	wire [6:0]fracture;
	
	Square uut(numberIn_tb, whole, fracture);
	
	initial begin
        numberIn_tb = 360;
        #5;
        numberIn_tb = 1;
        #5;
        numberIn_tb = 2;
        #5;
        numberIn_tb = 3;
        #5;
        numberIn_tb = 4;
        #5;
        numberIn_tb = 5;
        #5;
        numberIn_tb = 6;
        #5;
        numberIn_tb = 7;
        #5;
        numberIn_tb = 8;
        #5;
        numberIn_tb = 9;
        #5;
        numberIn_tb = 10;
        #5;
        numberIn_tb = 11;
        #5;
        numberIn_tb = 12;
        #5;
        numberIn_tb = 13;
        #5;
        numberIn_tb = 14;
        #5;
        numberIn_tb = 15;
        #5;
        numberIn_tb = 16;
        #5;
        numberIn_tb = 17;
        #5;
        numberIn_tb = 18;
        #5;
        numberIn_tb = 19;
        #5;
        numberIn_tb = 20;
        #5;
        numberIn_tb = 21;
        #5;
        numberIn_tb = 22;
        #5;
        numberIn_tb = 23;
        #5;
        numberIn_tb = 24;
        #5;
        numberIn_tb = 25;
        #5;
        numberIn_tb = 26;
        #5;
        numberIn_tb = 27;
        #5;
        numberIn_tb = 28;
        #5;
        numberIn_tb = 29;
        #5;
        numberIn_tb = 30;
        #5;
        numberIn_tb = 31;
        #5;
        numberIn_tb = 32;
        #5;
        numberIn_tb = 33;
        #5;
        numberIn_tb = 34;
        #5;
        numberIn_tb = 35;
        #5;
        numberIn_tb = 36;
        #5;
        numberIn_tb = 37;
        #5;
        numberIn_tb = 38;
        #5;
        numberIn_tb = 39;
        #5;
        numberIn_tb = 40;
        #5;
        numberIn_tb = 41;
        #5;
        numberIn_tb = 42;
        #5;
        numberIn_tb = 43;
        #5;
        numberIn_tb = 44;
        #5;
        numberIn_tb = 45;
        #5;
        numberIn_tb = 46;
        #5;
        numberIn_tb = 47;
        #5;
        numberIn_tb = 48;
        #5;
        numberIn_tb = 49;
        #5;
        numberIn_tb = 50;
        #5;
        numberIn_tb = 51;
        #5;
        numberIn_tb = 52;
        #5;
        numberIn_tb = 53;
        #5;
        numberIn_tb = 54;
        #5;
        numberIn_tb = 55;
        #5;
        numberIn_tb = 56;
        #5;
        numberIn_tb = 57;
        #5;
        numberIn_tb = 58;
        #5;
        numberIn_tb = 59;
        #5;
        numberIn_tb = 60;
        #5;
        numberIn_tb = 61;
        #5;
        numberIn_tb = 62;
        #5;
        numberIn_tb = 63;
        #5;
        numberIn_tb = 64;
        #5;
        numberIn_tb = 65;
        #5;
        numberIn_tb = 66;
        #5;
        numberIn_tb = 67;
        #5;
        numberIn_tb = 68;
        #5;
        numberIn_tb = 69;
        #5;
        numberIn_tb = 70;
        #5;
        numberIn_tb = 71;
        #5;
        numberIn_tb = 72;
        #5;
        numberIn_tb = 73;
        #5;
        numberIn_tb = 74;
        #5;
        numberIn_tb = 75;
        #5;
        numberIn_tb = 76;
        #5;
        numberIn_tb = 77;
        #5;
        numberIn_tb = 78;
        #5;
        numberIn_tb = 79;
        #5;
        numberIn_tb = 80;
        #5;
        numberIn_tb = 81;
        #5;
        numberIn_tb = 82;
        #5;
        numberIn_tb = 83;
        #5;
        numberIn_tb = 84;
        #5;
        numberIn_tb = 85;
        #5;
        numberIn_tb = 86;
        #5;
        numberIn_tb = 87;
        #5;
        numberIn_tb = 88;
        #5;
        numberIn_tb = 89;
        #5;
        numberIn_tb = 90;
        #5;
        numberIn_tb = 91;
        #5;
        numberIn_tb = 92;
        #5;
        numberIn_tb = 93;
        #5;
        numberIn_tb = 94;
        #5;
        numberIn_tb = 95;
        #5;
        numberIn_tb = 96;
        #5;
        numberIn_tb = 97;
        #5;
        numberIn_tb = 98;
        #5;
        numberIn_tb = 99;
        #5;
	end
	
endmodule
